library verilog;
use verilog.vl_types.all;
entity RCA8_vlg_vec_tst is
end RCA8_vlg_vec_tst;
